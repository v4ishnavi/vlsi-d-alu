magic
tech scmos
timestamp 1700598345
<< nwell >>
rect -26 6 48 28
rect 54 6 83 28
<< ntransistor >>
rect -14 -10 -12 -6
rect 2 -10 4 -6
rect 18 -10 20 -6
rect 34 -10 36 -6
rect 66 -11 68 -6
<< ptransistor >>
rect -14 12 -12 20
rect 2 12 4 20
rect 18 12 20 20
rect 34 12 36 20
rect 66 12 68 20
<< ndiffusion >>
rect -15 -10 -14 -6
rect -12 -10 -11 -6
rect 1 -10 2 -6
rect 4 -10 5 -6
rect 17 -10 18 -6
rect 20 -10 21 -6
rect 33 -10 34 -6
rect 36 -10 37 -6
rect 61 -7 66 -6
rect 65 -11 66 -7
rect 68 -10 69 -6
rect 68 -11 73 -10
<< pdiffusion >>
rect -15 16 -14 20
rect -19 12 -14 16
rect -12 12 2 20
rect 4 12 18 20
rect 20 12 34 20
rect 36 16 41 20
rect 36 12 37 16
rect 61 19 66 20
rect 65 15 66 19
rect 61 12 66 15
rect 68 16 73 20
rect 68 12 69 16
<< ndcontact >>
rect -19 -10 -15 -6
rect -11 -10 -7 -6
rect -3 -10 1 -6
rect 5 -10 9 -6
rect 13 -10 17 -6
rect 21 -10 25 -6
rect 29 -10 33 -6
rect 37 -10 41 -6
rect 61 -11 65 -7
rect 69 -10 73 -6
<< pdcontact >>
rect -19 16 -15 20
rect 37 12 41 16
rect 61 15 65 19
rect 69 12 73 16
<< polysilicon >>
rect -14 20 -12 34
rect 2 20 4 34
rect 18 20 20 34
rect 34 20 36 34
rect 66 20 68 23
rect -14 -6 -12 12
rect 2 -6 4 12
rect 18 -6 20 12
rect 34 -6 36 12
rect 66 3 68 12
rect 67 -1 68 3
rect 66 -6 68 -1
rect -14 -14 -12 -10
rect 2 -14 4 -10
rect 18 -14 20 -10
rect 34 -14 36 -10
rect 66 -14 68 -11
<< polycontact >>
rect -15 34 -11 38
rect 1 34 5 38
rect 17 34 21 38
rect 33 34 37 38
rect 63 -1 67 3
<< metal1 >>
rect -15 38 -10 41
rect -11 34 -10 38
rect 1 38 6 41
rect 5 34 6 38
rect 17 38 22 41
rect 21 34 22 38
rect 33 38 38 41
rect 37 34 38 38
rect -26 25 83 28
rect -18 20 -15 25
rect 62 19 65 25
rect 38 3 41 12
rect 70 3 73 12
rect -18 -1 63 3
rect 70 -1 81 3
rect -10 -6 -7 -1
rect 6 -6 9 -1
rect 22 -6 25 -1
rect 38 -6 41 -1
rect 70 -6 73 -1
rect -18 -16 -15 -10
rect -2 -16 1 -10
rect 14 -16 17 -10
rect 30 -16 33 -10
rect 62 -16 65 -11
rect -18 -20 67 -16
<< end >>
