magic
tech scmos
timestamp 1700473259
<< nwell >>
rect -39 8 -17 36
rect -8 8 16 36
rect 24 8 48 36
rect -8 -27 16 1
rect 24 -27 48 1
rect -39 -58 -17 -30
<< ntransistor >>
rect -32 -5 -28 -3
rect -1 -43 3 -41
rect 31 -42 35 -40
rect -1 -69 3 -67
rect 31 -69 35 -67
rect -32 -71 -28 -69
<< ptransistor >>
rect -32 21 -24 23
rect 0 21 8 23
rect 31 21 39 23
rect -1 -15 7 -13
rect 31 -15 39 -13
rect -32 -45 -24 -43
<< ndiffusion >>
rect -32 -3 -28 -2
rect -32 -7 -28 -5
rect -1 -36 3 -35
rect -1 -41 3 -40
rect -1 -44 3 -43
rect -1 -67 3 -65
rect 31 -40 35 -38
rect 31 -44 35 -42
rect 31 -67 35 -65
rect -32 -69 -28 -68
rect -32 -73 -28 -71
rect -1 -71 3 -69
rect 31 -71 35 -69
<< pdiffusion >>
rect -28 24 -24 28
rect -32 23 -24 24
rect 0 24 1 28
rect 5 24 8 28
rect 0 23 8 24
rect 31 24 32 28
rect 36 24 39 28
rect 31 23 39 24
rect -32 20 -24 21
rect -28 16 -24 20
rect 0 20 8 21
rect 0 16 1 20
rect 5 16 8 20
rect 31 20 39 21
rect 35 16 39 20
rect -1 -12 1 -8
rect 5 -12 7 -8
rect -1 -13 7 -12
rect 35 -12 39 -8
rect 31 -13 39 -12
rect -1 -16 7 -15
rect 3 -20 7 -16
rect -28 -42 -24 -38
rect -32 -43 -24 -42
rect -32 -46 -24 -45
rect -28 -50 -24 -46
rect 31 -16 39 -15
rect 35 -20 39 -16
<< ndcontact >>
rect -32 -2 -28 2
rect -32 -11 -28 -7
rect -1 -40 3 -36
rect -1 -48 3 -44
rect -32 -68 -28 -64
rect -1 -65 3 -61
rect 31 -38 35 -34
rect 31 -48 35 -44
rect 31 -65 35 -61
rect -32 -77 -28 -73
rect -1 -75 3 -71
rect 31 -75 35 -71
<< pdcontact >>
rect -32 24 -28 28
rect 1 24 5 28
rect 32 24 36 28
rect -32 16 -28 20
rect 1 16 5 20
rect 31 16 35 20
rect 1 -12 5 -8
rect 31 -12 35 -8
rect -1 -20 3 -16
rect -32 -42 -28 -38
rect -32 -50 -28 -46
rect 31 -20 35 -16
<< polysilicon >>
rect -57 39 -5 41
rect -57 10 -55 39
rect -7 23 -5 39
rect -44 21 -32 23
rect -24 21 -21 23
rect -7 21 0 23
rect 8 21 18 23
rect 22 21 31 23
rect 39 21 66 23
rect -44 10 -42 21
rect -57 8 -42 10
rect -57 -33 -55 8
rect -44 -3 -42 8
rect -44 -5 -32 -3
rect -28 -5 -24 -3
rect -44 -7 -42 -5
rect -6 -15 -1 -13
rect 7 -15 17 -13
rect 20 -15 31 -13
rect 39 -15 49 -13
rect -57 -35 -12 -33
rect -14 -41 -12 -35
rect -14 -43 -1 -41
rect 3 -43 6 -41
rect -44 -45 -32 -43
rect -24 -45 -21 -43
rect -44 -56 -42 -45
rect -50 -58 -42 -56
rect -87 -61 -64 -59
rect -87 -89 -85 -61
rect -50 -78 -48 -58
rect -44 -69 -42 -58
rect 20 -67 22 -15
rect 28 -42 31 -40
rect 35 -42 66 -40
rect -5 -69 -1 -67
rect 3 -69 22 -67
rect 28 -69 31 -67
rect 35 -69 45 -67
rect -44 -71 -32 -69
rect -28 -71 -24 -69
rect -44 -73 -42 -71
rect -5 -78 -3 -69
rect -50 -80 -3 -78
rect 43 -89 45 -69
rect -87 -91 45 -89
<< polycontact >>
rect 66 20 70 24
rect -10 -16 -6 -12
rect -64 -62 -60 -58
rect 66 -42 70 -38
<< metal1 >>
rect -49 44 75 47
rect -49 8 -46 44
rect -39 33 64 36
rect -31 28 -28 33
rect -31 8 -28 16
rect -49 5 -28 8
rect -31 2 -28 5
rect -31 -18 -28 -11
rect -77 -22 -28 -18
rect -77 -83 -74 -22
rect -16 -27 -13 33
rect 2 28 5 33
rect 33 28 36 33
rect 67 24 70 44
rect 2 -8 5 16
rect 32 -8 35 16
rect -31 -30 -13 -27
rect -31 -38 -28 -30
rect -31 -58 -28 -50
rect -60 -60 -28 -58
rect -10 -60 -7 -16
rect -1 -30 2 -20
rect 31 -30 34 -20
rect -1 -33 34 -30
rect -1 -36 2 -33
rect 31 -34 34 -33
rect 67 -38 70 20
rect 67 -43 70 -42
rect -60 -61 -7 -60
rect -31 -63 -7 -61
rect -1 -61 2 -48
rect 31 -61 34 -48
rect -31 -64 -28 -63
rect -31 -83 -28 -77
rect -1 -83 2 -75
rect 31 -83 34 -75
rect -77 -87 37 -83
rect -31 -88 -28 -87
rect -1 -88 2 -87
rect 31 -88 34 -87
<< end >>
