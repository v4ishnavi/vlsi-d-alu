magic
tech scmos
timestamp 1701334167
<< polysilicon >>
rect -275 257 562 259
rect -272 244 -270 257
rect 560 239 562 257
rect -219 233 331 235
rect 329 215 331 233
rect 329 213 341 215
rect -223 109 257 111
rect -223 -19 225 -17
rect -225 -140 196 -138
rect 19 -243 51 -241
rect -219 -281 -102 -279
rect -101 -351 -94 -349
rect 47 -382 51 -243
rect 2 -384 51 -382
rect -223 -405 -118 -403
rect -156 -406 -118 -405
rect -120 -486 -112 -484
rect 30 -525 33 -384
rect -1 -527 33 -525
rect -223 -533 -121 -531
rect -118 -633 -113 -630
rect -225 -654 -168 -652
rect -170 -680 -168 -654
rect 30 -669 33 -527
rect -14 -671 33 -669
rect -170 -684 -135 -680
rect 194 -738 196 -140
rect 223 -421 225 -19
rect 255 -97 257 109
rect 255 -99 328 -97
rect 784 -214 786 -213
rect 780 -216 786 -214
rect 285 -421 318 -419
rect 223 -423 287 -421
rect 194 -740 311 -738
rect -131 -750 -122 -748
<< polycontact >>
rect -273 239 -267 244
rect 547 239 551 243
rect 341 213 345 217
rect 13 -245 19 -239
rect -105 -351 -101 -347
rect -2 -385 2 -381
rect -124 -487 -120 -483
rect -5 -528 -1 -524
rect -124 -634 -118 -628
rect -18 -672 -14 -668
rect 547 -77 552 -72
rect 566 -77 570 -72
rect 328 -101 333 -96
rect 784 -213 788 -209
rect 547 -398 551 -394
rect 560 -396 564 -392
rect 318 -422 322 -418
rect 764 -539 768 -535
rect 548 -720 552 -716
rect 311 -741 315 -737
rect -136 -752 -131 -746
rect 755 -859 759 -855
<< metal1 >>
rect -325 259 -297 262
rect -301 256 -297 259
rect -301 252 -291 256
rect -301 156 -297 252
rect -272 232 -269 239
rect 548 236 551 239
rect 345 213 355 216
rect -187 72 337 77
rect -301 -357 -297 -236
rect -279 -252 -278 -247
rect -279 -282 -276 -252
rect -237 -282 -234 -240
rect -187 -256 -182 72
rect 548 -72 551 -60
rect 567 -85 570 -77
rect 333 -101 351 -97
rect 211 -158 342 -155
rect -184 -258 -182 -256
rect -279 -285 -272 -282
rect -237 -285 -227 -282
rect -110 -351 -105 -348
rect -227 -359 -122 -355
rect 211 -470 214 -158
rect 783 -209 786 -200
rect 783 -213 784 -209
rect 759 -363 764 -359
rect 769 -363 772 -361
rect 548 -394 551 -389
rect 561 -400 564 -396
rect 322 -422 350 -418
rect 82 -473 214 -470
rect 303 -479 339 -476
rect -128 -486 -124 -483
rect -232 -496 -136 -493
rect -232 -497 -230 -496
rect -225 -497 -136 -496
rect -287 -589 -286 -585
rect 303 -613 306 -479
rect 765 -535 768 -530
rect 83 -616 306 -613
rect -127 -633 -124 -629
rect -234 -640 -138 -636
rect 548 -716 551 -713
rect -237 -725 -153 -721
rect 315 -741 347 -738
rect 313 -743 347 -741
rect -141 -750 -136 -746
rect -279 -772 -276 -761
rect -327 -775 -276 -772
rect -241 -785 -237 -753
rect 82 -759 305 -756
rect -335 -789 -237 -785
rect -305 -803 -302 -789
rect 302 -797 305 -759
rect 302 -800 336 -797
rect -305 -806 -30 -803
rect -33 -894 -30 -806
rect 756 -855 759 -849
rect -33 -897 326 -894
rect 323 -1002 326 -897
rect 323 -1005 577 -1002
<< m2contact >>
rect 355 212 360 218
rect -287 178 -282 183
rect -290 55 -285 60
rect -291 -76 -286 -70
rect -294 -199 -289 -194
rect -278 -252 -273 -247
rect 337 71 343 77
rect 351 -102 356 -96
rect -85 -244 -80 -239
rect -189 -262 -184 -256
rect -35 -310 -30 -305
rect -288 -335 -283 -330
rect -115 -351 -110 -346
rect -52 -451 -47 -446
rect -290 -460 -285 -454
rect 77 -475 82 -469
rect 342 -160 348 -154
rect 350 -423 355 -417
rect -133 -487 -128 -482
rect -55 -594 -50 -589
rect 78 -617 83 -612
rect 339 -480 344 -475
rect -135 -634 -127 -627
rect -294 -714 -289 -708
rect -70 -739 -65 -734
rect 347 -743 353 -738
rect -148 -752 -141 -745
rect 77 -760 82 -755
rect 336 -801 341 -796
<< pdm12contact >>
rect -292 -590 -287 -584
<< metal2 >>
rect -314 179 -287 183
rect 331 156 353 159
rect 64 155 67 156
rect 331 155 334 156
rect 64 152 334 155
rect -319 55 -290 59
rect -318 -75 -291 -71
rect -318 -199 -294 -195
rect -214 -243 -85 -240
rect -214 -247 -210 -243
rect -273 -250 -210 -247
rect -326 -260 -189 -257
rect -184 -260 -177 -257
rect -315 -335 -288 -331
rect -180 -348 -177 -260
rect -34 -328 -31 -310
rect 64 -328 67 152
rect 758 133 949 137
rect 343 71 356 77
rect 801 61 842 64
rect 839 -65 842 61
rect 301 -68 842 -65
rect 301 -238 304 -68
rect 758 -181 921 -177
rect 301 -241 352 -238
rect 336 -243 352 -241
rect 797 -253 845 -250
rect -34 -331 67 -328
rect -180 -351 -115 -348
rect -314 -459 -290 -455
rect -180 -483 -177 -351
rect 842 -367 845 -253
rect 295 -370 845 -367
rect -51 -470 -48 -451
rect -51 -473 77 -470
rect -180 -486 -133 -483
rect -314 -589 -292 -585
rect -180 -629 -177 -486
rect 295 -558 298 -370
rect 753 -502 941 -498
rect 295 -561 350 -558
rect 796 -574 847 -571
rect -54 -613 -51 -594
rect -54 -616 78 -613
rect -180 -633 -135 -629
rect -320 -713 -294 -709
rect -180 -746 -177 -633
rect 844 -689 847 -574
rect 292 -692 847 -689
rect -180 -750 -148 -746
rect -69 -756 -66 -739
rect -69 -759 77 -756
rect 292 -880 295 -692
rect 750 -823 957 -819
rect 292 -883 348 -880
rect 793 -895 968 -892
<< m123contact >>
rect 547 231 552 236
rect 782 -52 787 -47
rect 547 -60 552 -55
rect 566 -90 571 -85
rect 782 -200 788 -195
rect 764 -363 769 -358
rect 547 -389 552 -384
rect 561 -405 566 -400
rect 764 -530 769 -525
rect 755 -685 760 -680
rect 547 -713 552 -708
rect 755 -849 760 -844
<< metal3 >>
rect 548 -55 551 231
rect 548 -89 566 -86
rect 548 -384 551 -89
rect 783 -195 786 -52
rect 548 -403 561 -400
rect 548 -708 551 -403
rect 765 -525 768 -363
rect 756 -844 759 -685
use enable  enable_1
timestamp 1700594004
transform 0 -1 -189 1 0 -632
box -129 30 358 112
use xor  xor_2
timestamp 1700473259
transform 1 0 -64 0 1 -560
box -87 -91 75 47
use xor  xor_3
timestamp 1700473259
transform 1 0 -78 0 1 -704
box -87 -91 75 47
use full_adder  full_adder_3
timestamp 1700594004
transform 1 0 533 0 1 -811
box -194 -197 263 108
use full_adder  full_adder_2
timestamp 1700594004
transform 1 0 536 0 1 -490
box -194 -197 263 108
use xor  xor_1
timestamp 1700473259
transform 1 0 -62 0 1 -417
box -87 -91 75 47
use enable  enable_0
timestamp 1700594004
transform 0 -1 -189 1 0 -118
box -129 30 358 112
use xor  xor_0
timestamp 1700473259
transform 1 0 -45 0 1 -276
box -87 -91 75 47
use full_adder  full_adder_0
timestamp 1700594004
transform 1 0 541 0 1 145
box -194 -197 263 108
use full_adder  full_adder_1
timestamp 1700594004
transform 1 0 537 0 1 -169
box -194 -197 263 108
<< end >>
