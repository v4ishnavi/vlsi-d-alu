magic
tech scmos
timestamp 1701329101
<< polysilicon >>
rect -94 484 -65 486
rect -98 360 -67 362
rect -98 232 -65 234
rect -33 189 181 190
rect 185 189 187 190
rect -33 188 187 189
rect -101 111 -63 113
rect -33 -16 -31 188
rect -94 -18 -31 -16
rect -3 77 -1 80
rect -3 75 184 77
rect -3 -140 -1 75
rect -99 -142 -1 -140
rect 42 -42 184 -40
rect 42 -268 44 -42
rect -99 -270 44 -268
rect 158 -169 185 -167
rect 158 -389 160 -169
rect -101 -391 160 -389
<< polycontact >>
rect -65 484 -61 488
rect -67 360 -63 364
rect -65 232 -61 236
rect 181 189 185 193
rect -63 111 -59 115
rect 184 75 188 79
rect 184 -42 188 -38
rect 185 -171 189 -167
<< metal1 >>
rect -100 501 246 504
rect -100 481 -97 501
rect -61 484 160 487
rect -242 432 -170 436
rect -174 404 -170 432
rect -63 360 148 363
rect -61 232 134 235
rect -59 111 124 114
rect -174 -101 -170 19
rect -152 -16 -149 5
rect -110 1 -107 15
rect -110 -2 -97 1
rect -152 -19 -142 -16
rect -145 -22 -142 -19
rect -100 -23 -97 -2
rect 121 -125 124 111
rect 131 -4 134 232
rect 145 115 148 360
rect 157 229 160 484
rect 243 275 246 501
rect 157 226 188 229
rect 185 189 188 192
rect 184 188 188 189
rect 198 172 201 178
rect 198 169 202 172
rect 199 163 202 169
rect 240 167 243 187
rect 240 164 247 167
rect 145 112 190 115
rect 188 75 189 78
rect 186 74 189 75
rect 199 47 202 63
rect 241 48 244 73
rect 199 45 203 47
rect 241 45 248 48
rect 199 44 202 45
rect 131 -7 191 -4
rect 188 -42 190 -41
rect 185 -45 190 -42
rect 200 -78 203 -56
rect 242 -75 245 -46
rect 242 -78 249 -75
rect 121 -128 193 -125
rect 186 -167 190 -164
rect 189 -168 190 -167
rect -161 -326 -159 -322
rect -153 -501 -148 -498
rect -151 -504 -148 -501
rect 200 -504 203 -179
rect -153 -507 203 -504
<< m2contact >>
rect 224 283 229 288
rect 225 169 230 174
rect 227 50 232 55
rect 227 -74 232 -69
<< metal2 >>
rect 229 283 248 286
rect 230 169 257 172
rect 232 50 264 53
rect 232 -73 264 -70
<< m123contact >>
rect -147 477 -142 482
rect -161 430 -156 435
rect -163 305 -158 311
rect -164 176 -159 181
rect -167 51 -162 57
rect -160 -73 -155 -67
rect -164 -196 -159 -191
rect -166 -326 -161 -321
rect -167 -450 -162 -445
rect -111 -492 -106 -487
<< metal3 >>
rect -168 477 -147 480
rect -184 430 -161 434
rect -184 429 -180 430
rect -242 425 -180 429
rect -251 306 -163 310
rect -255 176 -164 180
rect -254 52 -167 56
rect -252 -72 -160 -68
rect -259 -196 -164 -192
rect -260 -326 -166 -322
rect -258 -450 -167 -446
rect -110 -513 -107 -492
rect -262 -516 -107 -513
use and2  and2_3
timestamp 1700594004
transform 0 -1 217 1 0 -143
box -36 -31 73 27
use and2  and2_2
timestamp 1700594004
transform 0 -1 217 1 0 -20
box -36 -31 73 27
use and2  and2_1
timestamp 1700594004
transform 0 -1 216 1 0 99
box -36 -31 73 27
use and2  and2_0
timestamp 1700594004
transform 0 -1 215 1 0 213
box -36 -31 73 27
use enable  enable_1
timestamp 1700594004
transform 0 -1 -62 1 0 -369
box -129 30 358 112
use enable  enable_0
timestamp 1700594004
transform 0 -1 -62 1 0 133
box -129 30 358 112
<< end >>
