magic
tech scmos
timestamp 1700594004
<< nwell >>
rect -32 -8 -8 15
rect 5 -8 29 15
rect 41 -8 65 15
<< ntransistor >>
rect -21 -26 -19 -22
rect 16 -26 18 -22
rect 52 -26 54 -22
<< ptransistor >>
rect -21 -1 -19 7
rect 16 -1 18 7
rect 52 -1 54 7
<< ndiffusion >>
rect -22 -26 -21 -22
rect -19 -26 16 -22
rect 18 -26 52 -22
rect 54 -26 55 -22
<< pdiffusion >>
rect -22 3 -21 7
rect -26 -1 -21 3
rect -19 3 -14 7
rect -19 -1 -18 3
rect 15 3 16 7
rect 11 -1 16 3
rect 18 3 23 7
rect 18 -1 19 3
rect 51 3 52 7
rect 47 -1 52 3
rect 54 3 59 7
rect 54 -1 55 3
<< ndcontact >>
rect -26 -26 -22 -22
rect 55 -26 59 -22
<< pdcontact >>
rect -26 3 -22 7
rect -18 -1 -14 3
rect 11 3 15 7
rect 19 -1 23 3
rect 47 3 51 7
rect 55 -1 59 3
<< polysilicon >>
rect -21 7 -19 19
rect 16 7 18 19
rect 52 7 54 19
rect -21 -22 -19 -1
rect 16 -22 18 -1
rect 52 -22 54 -1
rect -21 -29 -19 -26
rect 16 -29 18 -26
rect 52 -29 54 -26
<< polycontact >>
rect -22 19 -18 23
rect 15 19 19 23
rect 51 19 55 23
<< metal1 >>
rect -22 23 -18 25
rect 15 23 19 25
rect 51 23 55 25
rect -32 12 73 15
rect -25 7 -22 12
rect 12 7 15 12
rect 48 7 51 12
rect -18 -11 -15 -1
rect 19 -11 22 -1
rect 55 -11 58 -1
rect -18 -12 63 -11
rect -18 -13 66 -12
rect -18 -15 73 -13
rect 56 -22 59 -15
rect 63 -17 73 -15
rect 97 -16 103 -13
rect -26 -32 -23 -26
rect 66 -32 74 -30
rect -26 -33 74 -32
rect -26 -35 69 -33
use not  not_0
timestamp 1700473189
transform 1 0 85 0 1 0
box -12 -33 12 15
<< end >>
