magic
tech scmos
timestamp 1700473189
<< nwell >>
rect -12 -9 12 15
<< ntransistor >>
rect -1 -25 1 -21
<< ptransistor >>
rect -1 -2 1 6
<< ndiffusion >>
rect -3 -25 -1 -21
rect 1 -25 2 -21
<< pdiffusion >>
rect -2 2 -1 6
rect -6 -2 -1 2
rect 1 2 2 6
rect 1 -2 6 2
<< ndcontact >>
rect -7 -25 -3 -21
rect 2 -25 6 -21
<< pdcontact >>
rect -6 2 -2 6
rect 2 2 6 6
<< polysilicon >>
rect -1 6 1 9
rect -1 -14 1 -2
rect -5 -16 1 -14
rect -1 -21 1 -16
rect -1 -28 1 -25
<< polycontact >>
rect -9 -17 -5 -13
<< metal1 >>
rect -12 12 12 15
rect -5 6 -2 12
rect 2 -13 5 2
rect -12 -17 -9 -13
rect 2 -16 12 -13
rect 2 -21 5 -16
rect -6 -30 -3 -25
rect -12 -33 12 -30
<< end >>
