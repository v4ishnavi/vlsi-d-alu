magic
tech scmos
timestamp 1700594004
<< polysilicon >>
rect -13 94 48 96
rect 46 81 48 94
rect 178 72 192 74
rect -21 -55 -19 -3
rect 188 -47 243 -45
rect -21 -57 85 -55
rect -21 -58 -19 -57
rect 83 -63 85 -57
rect 241 -100 243 -47
rect 136 -127 145 -125
rect 142 -192 145 -127
<< polycontact >>
rect -17 93 -13 97
rect 45 77 49 81
rect -136 68 -132 72
rect 174 71 178 75
rect 192 71 196 75
rect 54 46 58 50
rect -123 10 -119 14
rect -22 -3 -18 1
rect 61 -33 65 -29
rect 184 -48 188 -44
rect 82 -67 86 -63
rect 241 -104 245 -100
rect 132 -127 136 -123
rect 141 -196 145 -192
<< metal1 >>
rect 45 74 48 77
rect -146 68 -136 71
rect -178 -136 -174 10
rect -170 -130 -167 67
rect 47 46 54 49
rect -135 10 -123 13
rect -22 1 -19 9
rect -40 -26 16 -22
rect 12 -43 16 -26
rect 58 -32 61 -29
rect 12 -48 38 -43
rect 150 -48 184 -44
rect 82 -69 86 -67
rect 192 -79 196 71
rect 134 -82 199 -79
rect 196 -101 199 -82
rect -170 -133 86 -130
rect -178 -140 49 -136
rect 82 -140 86 -133
rect 132 -144 198 -141
rect 132 -149 135 -144
rect 196 -145 198 -144
rect 186 -152 187 -148
rect 135 -196 141 -194
rect 242 -194 245 -174
rect 145 -196 245 -194
rect 135 -197 245 -196
<< m2contact >>
rect -171 67 -166 72
rect -152 67 -146 73
rect 45 69 50 74
rect 73 70 78 75
rect -179 10 -174 15
rect 42 46 47 51
rect -66 27 -61 32
rect -141 9 -135 15
rect -24 9 -18 15
rect 122 4 128 10
rect 53 -33 58 -28
rect 44 -71 49 -66
rect 223 -93 228 -88
rect 139 -111 145 -105
rect 180 -153 186 -147
rect 180 -173 186 -167
rect 140 -182 147 -175
<< metal2 >>
rect -184 68 -171 72
rect -166 68 -152 72
rect 50 71 73 74
rect 15 46 42 49
rect -66 16 -63 27
rect 15 16 18 46
rect -66 15 18 16
rect -194 10 -179 14
rect -174 10 -141 14
rect -66 13 -24 15
rect -66 12 -63 13
rect -18 13 18 15
rect 123 -8 127 4
rect 123 -12 221 -8
rect 3 -33 53 -29
rect 3 -58 8 -33
rect 3 -62 49 -58
rect 3 -68 8 -62
rect 45 -66 49 -62
rect -187 -74 8 -68
rect 224 -84 263 -81
rect 224 -88 227 -84
rect 145 -110 176 -107
rect 172 -148 176 -110
rect 172 -152 180 -148
rect 179 -173 180 -168
rect 179 -177 183 -173
rect 147 -180 183 -177
use xor  xor_1
timestamp 1700473259
transform 1 0 114 0 1 39
box -87 -91 75 47
use xor  xor_0
timestamp 1700473259
transform 1 0 -76 0 1 61
box -87 -91 75 47
use and2  and2_0
timestamp 1700594004
transform 1 0 70 0 1 -96
box -36 -31 73 27
use and2  and2_1
timestamp 1700594004
transform 1 0 70 0 1 -166
box -36 -31 73 27
use or2  or2_0
timestamp 1700594004
transform 0 -1 228 1 0 -169
box -13 -17 76 42
<< end >>
