magic
tech scmos
timestamp 1700594004
<< nwell >>
rect -13 8 31 32
<< ntransistor >>
rect -2 -7 0 -3
rect 18 -7 20 -3
<< ptransistor >>
rect -2 16 0 24
rect 18 16 20 24
<< ndiffusion >>
rect -3 -7 -2 -3
rect 0 -7 1 -3
rect 17 -7 18 -3
rect 20 -7 21 -3
<< pdiffusion >>
rect -3 20 -2 24
rect -7 16 -2 20
rect 0 16 18 24
rect 20 20 25 24
rect 20 16 21 20
<< ndcontact >>
rect -7 -7 -3 -3
rect 1 -7 5 -3
rect 13 -7 17 -3
rect 21 -7 25 -3
<< pdcontact >>
rect -7 20 -3 24
rect 21 16 25 20
<< polysilicon >>
rect -2 24 0 35
rect 18 24 20 35
rect -2 -3 0 16
rect 18 -3 20 16
rect -2 -12 0 -7
rect 18 -12 20 -7
<< polycontact >>
rect -3 35 1 39
rect 17 35 21 39
<< metal1 >>
rect -3 39 1 42
rect 17 39 21 42
rect -13 29 45 32
rect -6 24 -3 29
rect 22 5 25 16
rect -7 4 47 5
rect -7 2 44 4
rect 2 -3 5 2
rect 22 -3 25 2
rect 68 1 76 4
rect -6 -14 -3 -7
rect 14 -14 17 -7
rect 41 -14 44 -13
rect -6 -17 44 -14
use not  not_0
timestamp 1700473189
transform 1 0 56 0 1 17
box -12 -33 12 15
<< end >>
