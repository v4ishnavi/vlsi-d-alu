magic
tech scmos
timestamp 1700594004
<< polysilicon >>
rect -307 117 -285 119
rect -313 -27 -288 -25
rect -112 -42 -47 -40
rect -304 -169 -294 -167
rect 4 -227 6 -216
rect -116 -229 6 -227
rect -323 -313 -305 -311
<< polycontact >>
rect -278 38 -274 42
rect -116 -42 -112 -38
rect -51 -46 -47 -42
rect -283 -105 -279 -101
rect 3 -216 7 -212
rect -120 -230 -116 -226
rect -287 -248 -283 -244
rect -298 -392 -294 -388
<< metal1 >>
rect -97 74 -90 77
rect -281 39 -278 42
rect -283 38 -278 39
rect -93 -61 -90 74
rect -21 -33 25 -30
rect -21 -37 -18 -33
rect -47 -46 -46 -43
rect -49 -50 -46 -46
rect -93 -64 -65 -61
rect -103 -70 -86 -67
rect -285 -105 -283 -102
rect -285 -106 -281 -105
rect -89 -135 -86 -70
rect -68 -96 -65 -64
rect -68 -99 -57 -96
rect -89 -138 -59 -135
rect -87 -174 -60 -171
rect -87 -209 -84 -174
rect -108 -212 -84 -209
rect -76 -211 -59 -208
rect -76 -216 -73 -211
rect -100 -219 -73 -216
rect -295 -245 -287 -244
rect -291 -247 -287 -245
rect -100 -353 -97 -219
rect -119 -356 -97 -353
rect -305 -389 -298 -388
rect -301 -391 -298 -389
<< m2contact >>
rect -286 39 -281 44
rect -290 -107 -285 -102
rect -296 -250 -291 -245
rect -306 -394 -301 -389
<< metal2 >>
rect -310 39 -286 41
rect -310 38 -281 39
rect -312 -106 -290 -103
rect -320 -245 -292 -244
rect -320 -247 -296 -245
rect -327 -389 -303 -388
rect -327 -391 -306 -389
<< m123contact >>
rect -256 141 -251 146
rect -166 141 -161 146
rect -293 22 -288 27
rect -174 -2 -169 3
rect -294 -57 -289 -52
rect -295 -123 -290 -118
rect -186 -143 -181 -138
rect -295 -199 -290 -194
rect -298 -266 -292 -261
rect -186 -288 -181 -283
rect -300 -342 -295 -337
rect -305 -408 -300 -403
<< metal3 >>
rect -303 142 -256 145
rect -293 -52 -290 22
rect -165 7 -162 141
rect -172 4 -162 7
rect -172 3 -164 4
rect -169 -2 -164 3
rect -294 -194 -291 -123
rect -167 -134 -164 -2
rect -184 -137 -164 -134
rect -184 -138 -181 -137
rect -297 -337 -293 -266
rect -175 -278 -172 -137
rect -184 -281 -172 -278
rect -184 -283 -181 -281
rect -295 -341 -293 -337
rect -304 -419 -300 -408
rect -358 -423 -300 -419
use xnor  xnor_0
timestamp 1700594004
transform 1 0 -98 0 1 51
box -205 -33 2 105
use xnor  xnor_1
timestamp 1700594004
transform 1 0 -103 0 1 -93
box -205 -33 2 105
use xnor  xnor_2
timestamp 1700594004
transform 1 0 -107 0 1 -235
box -205 -33 2 105
use xnor  xnor_3
timestamp 1700594004
transform 1 0 -118 0 1 -379
box -205 -33 2 105
use and4  and4_0
timestamp 1700594004
transform 0 -1 -26 1 0 -182
box -40 -32 146 34
<< end >>
