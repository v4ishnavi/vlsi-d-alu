magic
tech scmos
timestamp 1701341286
<< polysilicon >>
rect -371 1175 -340 1177
rect -1453 1000 -1208 1002
rect -1453 -350 -1451 1000
rect -1210 966 -1208 1000
rect -1287 964 -1007 966
rect -1291 840 -1198 842
rect -1194 840 -1031 842
rect -1291 712 -1244 714
rect -1240 712 -1168 714
rect -1164 712 -1078 714
rect -1293 591 -1280 593
rect -1276 591 -1106 593
rect -1286 227 -1284 229
rect -1108 146 -1106 591
rect -1080 290 -1078 712
rect -1033 432 -1031 840
rect -1009 746 -1007 964
rect -1009 744 -721 746
rect -1009 576 -1007 744
rect -723 726 -721 744
rect -1009 574 -928 576
rect -1009 572 -1007 574
rect -1033 430 -930 432
rect -1033 429 -1031 430
rect -597 424 -404 426
rect -1080 288 -922 290
rect -1108 144 -943 146
rect -1108 142 -1106 144
rect -1180 114 -1179 116
rect -1175 114 -1036 116
rect -1290 103 -1289 105
rect -1038 -313 -1036 114
rect -642 87 -640 89
rect -750 85 -640 87
rect -642 -5 -640 85
rect -379 -201 -346 -199
rect -1038 -315 -711 -313
rect -1453 -352 -844 -350
rect -846 -648 -844 -352
rect -713 -448 -711 -315
rect -713 -450 -673 -448
rect -713 -451 -711 -450
rect -846 -650 -793 -648
<< polycontact >>
rect -376 1174 -371 1179
rect -1198 839 -1194 843
rect -1244 711 -1240 715
rect -1168 712 -1164 716
rect -1280 590 -1276 594
rect -1284 226 -1280 230
rect -726 721 -721 726
rect -601 423 -597 428
rect -1179 113 -1175 117
rect -1289 102 -1285 106
rect -1289 -26 -1285 -22
rect -1292 -147 -1288 -143
rect -754 84 -750 88
rect -384 -202 -379 -198
rect -673 -451 -669 -447
rect -793 -650 -789 -646
<< metal1 >>
rect -1279 1335 -659 1338
rect -1279 990 -1276 1335
rect -662 1329 -659 1335
rect -1430 987 -1276 990
rect -1430 -264 -1427 987
rect -1354 910 -1351 914
rect -1393 891 -1364 895
rect -1398 146 -1394 889
rect -1368 888 -1364 891
rect -1354 786 -1353 790
rect -1354 656 -1351 660
rect -1279 594 -1276 987
rect -1257 1243 -686 1247
rect -1356 532 -1354 536
rect -1346 474 -1343 484
rect -1346 471 -1335 474
rect -1338 226 -1335 471
rect -1304 259 -1301 494
rect -1304 256 -1290 259
rect -1293 224 -1290 256
rect -1280 227 -1277 230
rect -1257 212 -1253 1243
rect -1243 1183 -681 1186
rect -1243 715 -1240 1183
rect -684 1177 -681 1183
rect -1221 1108 -684 1111
rect -1273 208 -1253 212
rect -1351 173 -1350 177
rect -1398 142 -1363 146
rect -1285 103 -1282 106
rect -1285 -25 -1282 -22
rect -1273 -142 -1269 208
rect -1221 0 -1218 1108
rect -970 1088 -685 1091
rect -1148 894 -1042 897
rect -1197 843 -1194 849
rect -1148 826 -1145 894
rect -1185 823 -1145 826
rect -1185 117 -1182 823
rect -1167 709 -1164 712
rect -970 636 -967 1088
rect -688 1074 -685 1088
rect -688 1071 -644 1074
rect -691 925 -638 928
rect -659 900 -638 903
rect -659 897 -656 900
rect -693 894 -656 897
rect -695 847 -665 850
rect -668 845 -665 847
rect -668 842 -637 845
rect -644 775 -641 792
rect -680 772 -641 775
rect -721 723 -639 726
rect -722 713 -663 716
rect -666 707 -663 713
rect -666 704 -639 707
rect -970 633 -548 636
rect -1185 114 -1179 117
rect -1185 108 -1182 114
rect -1221 -3 -1200 0
rect -1221 -21 -1218 -3
rect -1288 -146 -1284 -143
rect -1203 -171 -1200 -3
rect -1151 -157 -1148 226
rect -551 194 -548 633
rect -723 191 -548 194
rect -931 -124 -665 -121
rect -1203 -174 -965 -171
rect -931 -264 -928 -124
rect -668 -125 -665 -124
rect -668 -128 -655 -125
rect -1430 -267 -928 -264
rect -1430 -291 -1427 -267
rect -669 -451 -650 -448
rect -682 -475 -649 -473
rect -701 -476 -649 -475
rect -701 -478 -679 -476
rect -644 -476 -642 -473
rect -763 -532 -760 -513
rect -763 -535 -649 -532
rect -789 -649 -674 -647
rect -789 -650 -649 -649
rect -677 -652 -649 -650
rect -677 -654 -674 -652
<< m2contact >>
rect -663 1324 -658 1329
rect -686 1243 -681 1248
rect -1277 226 -1272 231
rect -685 1172 -680 1177
rect -1282 102 -1277 107
rect -1282 -26 -1277 -21
rect -684 1106 -678 1111
rect -1198 849 -1193 854
rect -1042 893 -1037 898
rect -1168 704 -1163 709
rect -644 1070 -639 1075
rect -696 925 -691 930
rect -638 924 -633 929
rect -638 899 -633 904
rect -700 847 -695 852
rect -637 841 -632 846
rect -644 792 -639 797
rect -685 771 -680 776
rect -639 722 -633 728
rect -727 712 -722 717
rect -639 704 -634 709
rect -700 318 -695 323
rect -701 283 -696 288
rect -1152 226 -1147 231
rect -1186 103 -1181 108
rect -1222 -26 -1217 -21
rect -1284 -147 -1279 -142
rect -1273 -147 -1268 -142
rect -965 -175 -960 -170
rect -655 -129 -650 -124
rect -650 -452 -644 -446
rect -706 -478 -701 -473
rect -649 -477 -644 -472
rect -649 -535 -644 -530
rect -649 -653 -644 -648
<< pdm12contact >>
rect -698 894 -693 899
<< metal2 >>
rect -658 1326 -635 1329
rect -677 1248 -637 1251
rect -677 1247 -674 1248
rect -681 1244 -674 1247
rect -680 1174 -634 1177
rect -678 1107 -635 1110
rect -1197 925 -696 928
rect -1197 876 -1194 925
rect -1037 894 -698 897
rect -1443 873 -1194 876
rect -1443 -327 -1440 873
rect -1197 854 -1194 873
rect -953 713 -727 716
rect -1167 700 -1164 704
rect -1418 697 -1164 700
rect -1418 -288 -1415 697
rect -1072 497 -1069 505
rect -953 497 -950 713
rect -722 713 -721 716
rect -934 497 -933 498
rect -1072 494 -931 497
rect -1272 227 -1152 230
rect -1072 230 -1069 494
rect -698 441 -695 847
rect -684 620 -681 771
rect -684 617 -556 620
rect -1147 227 -1069 230
rect -1032 351 -933 354
rect -1277 103 -1186 106
rect -1032 106 -1029 351
rect -698 323 -695 436
rect -1181 103 -1029 106
rect -1006 213 -1003 214
rect -1006 210 -941 213
rect -1277 -25 -1222 -22
rect -1006 -22 -1003 210
rect -699 205 -696 283
rect -559 205 -556 617
rect -699 202 -556 205
rect -670 102 -667 202
rect -714 99 -667 102
rect -1217 -25 -1003 -22
rect -977 69 -974 70
rect -977 66 -948 69
rect -977 -38 -974 66
rect -714 69 -711 99
rect -727 66 -711 69
rect -977 -41 -658 -38
rect -1279 -146 -1273 -143
rect -977 -143 -974 -41
rect -661 -47 -658 -41
rect -661 -50 -644 -47
rect -661 -51 -658 -50
rect -650 -128 -647 -125
rect -1268 -146 -974 -143
rect -960 -174 -647 -171
rect -650 -202 -647 -174
rect -913 -268 -910 -267
rect -655 -268 -644 -266
rect -913 -269 -644 -268
rect -913 -271 -652 -269
rect -913 -288 -910 -271
rect -1418 -291 -910 -288
rect -1443 -330 -721 -327
rect -724 -475 -721 -330
rect -724 -478 -706 -475
<< m3contact >>
rect -700 436 -695 441
rect -733 65 -727 71
rect -657 -295 -652 -290
rect -658 -583 -653 -578
rect -637 -673 -632 -668
<< m123contact >>
rect -1341 954 -1336 959
rect -566 955 -561 960
rect -1359 909 -1354 915
rect -1399 889 -1393 896
rect -1360 785 -1354 791
rect -1359 656 -1354 661
rect -1302 648 -1297 653
rect -1347 598 -1342 603
rect -1361 531 -1356 536
rect -521 652 -516 657
rect -1357 172 -1351 178
rect -1357 49 -1352 54
rect -1299 33 -1294 38
rect -758 129 -753 134
rect -731 100 -726 105
rect -1357 -81 -1352 -76
rect -577 -140 -572 -135
rect -1152 -162 -1147 -157
rect -1360 -206 -1355 -201
rect -1304 -247 -1299 -242
rect -1346 -254 -1341 -249
rect -764 -513 -759 -508
<< metal3 >>
rect -1336 955 -566 958
rect -1507 910 -1359 914
rect -1510 891 -1399 895
rect -1513 786 -1360 790
rect -1526 656 -1359 660
rect -1297 649 -518 652
rect -1342 599 -924 602
rect -1531 532 -1361 536
rect -695 437 -535 440
rect -1530 173 -1357 177
rect -753 130 -605 133
rect -729 87 -726 100
rect -729 84 -674 87
rect -731 61 -728 65
rect -731 58 -687 61
rect -1526 49 -1357 53
rect -1300 34 -1299 38
rect -1294 34 -979 38
rect -1525 -81 -1357 -77
rect -1528 -205 -1360 -201
rect -1521 -253 -1346 -250
rect -1303 -268 -1300 -247
rect -1518 -271 -1300 -268
rect -1151 -509 -1148 -162
rect -1151 -512 -764 -509
rect -690 -601 -687 58
rect -677 -291 -674 84
rect -608 -135 -605 130
rect -538 16 -535 437
rect -538 13 -387 16
rect -608 -136 -581 -135
rect -608 -138 -577 -136
rect -584 -139 -577 -138
rect -677 -294 -657 -291
rect -390 -335 -387 13
rect -477 -338 -387 -335
rect -657 -601 -654 -583
rect -690 -604 -654 -601
rect -636 -753 -633 -673
rect -477 -753 -474 -338
rect -636 -756 -474 -753
use comparator  comparator_1
timestamp 1700600503
transform 0 1 -549 -1 0 -396
box -401 -116 331 166
use comparator  comparator_0
timestamp 1700600503
transform 0 1 -538 -1 0 980
box -401 -116 331 166
use equal  equal_0
timestamp 1700594004
transform 1 0 -623 0 1 457
box -358 -423 25 156
use enable  enable_1
timestamp 1700594004
transform 0 -1 -1255 1 0 -124
box -129 30 358 112
use enable  enable_0
timestamp 1700594004
transform 0 -1 -1256 1 0 613
box -129 30 358 112
<< end >>
