magic
tech scmos
timestamp 1700600503
<< nwell >>
rect -181 -77 -157 -53
rect -3 -74 21 -50
rect 198 -78 222 -54
<< ntransistor >>
rect 33 -63 37 -61
rect -145 -66 -141 -64
rect 234 -67 238 -65
<< ptransistor >>
rect 6 -63 14 -61
rect -172 -66 -164 -64
rect 207 -67 215 -65
<< ndiffusion >>
rect 33 -61 37 -60
rect -145 -64 -141 -63
rect -145 -68 -141 -66
rect 33 -65 37 -63
rect 234 -65 238 -64
rect 234 -69 238 -67
<< pdiffusion >>
rect -168 -63 -164 -59
rect -172 -64 -164 -63
rect 10 -60 14 -56
rect 6 -61 14 -60
rect 6 -64 14 -63
rect -172 -67 -164 -66
rect -168 -71 -164 -67
rect 10 -68 14 -64
rect 211 -64 215 -60
rect 207 -65 215 -64
rect 207 -68 215 -67
rect 211 -72 215 -68
<< ndcontact >>
rect -145 -63 -141 -59
rect 33 -60 37 -56
rect -145 -72 -141 -68
rect 33 -69 37 -65
rect 234 -64 238 -60
rect 234 -73 238 -69
<< pdcontact >>
rect -172 -63 -168 -59
rect 6 -60 10 -56
rect -172 -71 -168 -67
rect 6 -68 10 -64
rect 207 -64 211 -60
rect 207 -72 211 -68
<< polysilicon >>
rect -351 142 -182 144
rect -351 115 -349 142
rect -392 113 -349 115
rect -392 -95 -390 113
rect -351 24 -349 113
rect -94 36 -92 38
rect 117 36 119 41
rect -375 4 -372 23
rect -351 19 -349 20
rect -246 4 -244 27
rect -94 4 -92 32
rect 117 4 119 32
rect -283 -61 -269 -60
rect -283 -62 -272 -61
rect 3 -63 6 -61
rect 14 -63 33 -61
rect 37 -62 54 -61
rect 37 -63 52 -62
rect -175 -66 -172 -64
rect -164 -66 -145 -64
rect -141 -66 -128 -64
rect -152 -70 -150 -66
rect -280 -90 -278 -72
rect 26 -67 28 -63
rect 204 -67 207 -65
rect 215 -67 234 -65
rect 238 -67 256 -65
rect 227 -71 229 -67
rect 42 -73 44 -72
rect -136 -75 -134 -74
rect 254 -68 256 -67
rect -136 -90 -134 -79
rect 42 -90 44 -77
rect 243 -90 245 -79
rect -280 -92 245 -90
rect -260 -95 -258 -92
rect -392 -97 -258 -95
rect -260 -99 -258 -97
<< polycontact >>
rect -182 142 -178 146
rect -375 23 -370 29
rect -94 32 -90 36
rect 116 32 120 36
rect -247 27 -243 31
rect -352 20 -348 24
rect -376 0 -372 4
rect -248 0 -244 4
rect -96 0 -92 4
rect 115 0 119 4
rect -272 -65 -268 -61
rect -281 -72 -277 -68
rect -153 -74 -149 -70
rect -130 -70 -126 -66
rect 25 -71 29 -67
rect 52 -66 56 -62
rect -137 -79 -133 -75
rect 41 -77 45 -73
rect 226 -75 230 -71
rect 254 -72 258 -68
rect 242 -79 246 -75
<< metal1 >>
rect -198 121 -194 166
rect -401 96 -197 99
rect -401 -25 -398 96
rect -152 81 -149 84
rect -375 78 -149 81
rect -375 29 -372 78
rect -136 50 -133 83
rect -247 47 -133 50
rect -247 31 -244 47
rect -118 44 -115 84
rect -104 53 -101 86
rect -104 50 119 53
rect -118 41 -91 44
rect -118 38 -115 41
rect -94 36 -91 41
rect 116 36 119 50
rect 84 21 131 24
rect -276 18 -239 21
rect -119 18 -86 21
rect -369 -25 -367 -24
rect -401 -28 -366 -25
rect -307 -26 -304 -25
rect -309 -27 -304 -26
rect -268 -27 -237 -24
rect -112 -27 -86 -24
rect 90 -27 123 -24
rect -318 -38 -315 -35
rect -349 -41 -315 -38
rect -349 -44 -346 -41
rect -307 -44 -304 -27
rect -326 -47 -304 -44
rect -298 -40 -277 -37
rect -326 -51 -323 -47
rect -298 -52 -295 -40
rect -197 -44 -194 -35
rect -125 -37 -121 -35
rect -162 -40 -150 -37
rect -271 -67 -268 -65
rect -181 -67 -178 -53
rect -153 -60 -150 -40
rect -168 -63 -145 -60
rect -181 -70 -172 -67
rect -326 -76 -323 -73
rect -181 -76 -178 -70
rect -136 -68 -133 -53
rect -125 -56 -122 -37
rect -34 -55 -31 -36
rect 4 -40 7 -36
rect -21 -43 7 -40
rect 25 -41 44 -38
rect -21 -53 -18 -43
rect -125 -59 -106 -56
rect -109 -62 -106 -59
rect -326 -79 -178 -76
rect -141 -71 -133 -68
rect -153 -77 -149 -74
rect -136 -75 -133 -71
rect -109 -68 -106 -67
rect -3 -64 0 -50
rect 25 -57 28 -41
rect 77 -47 81 -37
rect 135 -43 170 -39
rect 135 -44 139 -43
rect 10 -60 33 -57
rect -3 -67 6 -64
rect -130 -73 -127 -70
rect -181 -83 -178 -79
rect -3 -83 0 -67
rect 42 -65 45 -50
rect 182 -44 208 -40
rect 241 -41 257 -37
rect 182 -47 186 -44
rect 279 -47 282 -40
rect 316 -42 320 -38
rect 317 -46 320 -42
rect 185 -52 186 -47
rect 226 -50 282 -47
rect 37 -68 45 -65
rect 25 -74 29 -71
rect 42 -73 45 -68
rect 52 -69 55 -66
rect 198 -68 201 -54
rect 226 -61 229 -50
rect 211 -64 234 -61
rect 198 -71 207 -68
rect 198 -83 201 -71
rect 243 -69 246 -54
rect 238 -72 246 -69
rect 243 -75 246 -72
rect 226 -78 230 -75
rect 254 -75 257 -72
rect -181 -86 201 -83
<< m2contact >>
rect -350 -49 -345 -44
rect -199 -49 -194 -44
rect -271 -72 -266 -67
rect -35 -60 -30 -55
rect -22 -58 -17 -53
rect -111 -67 -106 -62
rect -130 -78 -125 -73
rect 76 -52 81 -47
rect 133 -50 139 -44
rect 257 -41 263 -36
rect 180 -52 185 -47
rect 316 -51 321 -46
rect 52 -74 57 -69
rect 254 -81 260 -75
<< metal2 >>
rect -349 -44 -346 -43
rect -349 -99 -346 -49
rect -271 -99 -268 -72
rect -197 -99 -194 -49
rect -130 -97 -127 -78
rect -109 -102 -106 -67
rect -34 -102 -31 -60
rect -109 -105 -31 -102
rect -34 -113 -31 -105
rect -21 -105 -18 -58
rect 52 -98 55 -74
rect 77 -97 81 -52
rect 135 -97 139 -50
rect 182 -105 185 -52
rect 258 -54 262 -41
rect 258 -58 276 -54
rect 254 -99 257 -81
rect 272 -98 276 -58
rect -21 -108 185 -105
rect 317 -113 320 -51
rect -34 -116 322 -113
use and5  and5_0
timestamp 1700594041
transform -1 0 319 0 -1 -17
box -12 -41 202 24
use and4  and4_0
timestamp 1700594004
transform -1 0 52 0 -1 -4
box -40 -32 146 34
use and3  and3_0
timestamp 1700594004
transform -1 0 -143 0 -1 -12
box -32 -35 103 25
use and2  and2_0
timestamp 1700594004
transform -1 0 -302 0 -1 -10
box -36 -31 73 27
use not  not_0
timestamp 1700473189
transform 0 -1 -311 1 0 -61
box -12 -33 12 15
use or4  or4_0
timestamp 1700598345
transform -1 0 -114 0 -1 124
box -26 -20 83 41
<< end >>
