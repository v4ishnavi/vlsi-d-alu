magic
tech scmos
timestamp 1701520041
<< polysilicon >>
rect 2197 1724 2278 1726
rect 15 1309 23 1311
rect 15 243 17 1309
rect 28 1309 42 1311
rect 2218 1054 2324 1056
rect 2218 1035 2220 1054
rect 2133 973 2169 975
rect 2127 940 2129 942
rect 2127 938 2172 940
rect 2127 892 2129 938
rect 2127 890 2389 892
rect 2190 348 2219 350
rect -279 241 17 243
rect -281 120 -222 122
rect -644 74 -435 76
rect -422 54 -416 56
rect -281 6 -248 8
rect -224 -6 -222 120
rect 583 92 1292 94
rect -224 -8 -46 -6
rect -224 -84 -222 -8
rect -224 -86 -160 -84
rect -276 -104 -154 -102
rect -48 -727 -46 -8
rect 1290 -145 1292 92
rect 1290 -147 1771 -145
rect 1769 -265 1771 -147
rect 2387 -265 2389 890
rect 1769 -267 2389 -265
rect -48 -729 293 -727
<< polycontact >>
rect 23 1308 28 1313
rect 2217 1031 2221 1035
rect 2169 972 2173 976
rect 2172 936 2176 941
rect -426 53 -422 57
rect -248 6 -244 10
rect 579 91 583 95
rect -160 -87 -156 -83
rect -154 -105 -150 -100
rect 1011 -215 1016 -211
rect 293 -729 297 -725
<< metal1 >>
rect 2022 1219 2237 1222
rect 1974 1191 1977 1200
rect 1972 1188 2192 1191
rect 2189 1023 2192 1188
rect 2234 1024 2237 1219
rect 2170 976 2180 978
rect 2173 974 2180 976
rect 2176 937 2180 941
rect 1012 296 1016 299
rect -137 94 -50 97
rect -644 54 -426 57
rect -137 9 -134 94
rect -45 94 -25 97
rect 574 95 582 96
rect 574 92 579 95
rect -244 6 -134 9
rect -97 -15 -7 -12
rect -97 -30 -94 -15
rect -138 -81 -134 -80
rect -138 -84 -135 -81
rect -156 -87 -135 -84
rect -150 -104 -135 -101
rect -79 -122 -76 -104
rect -288 -125 -76 -122
rect -156 -151 -153 -140
rect -156 -154 -71 -151
rect -292 -1254 -288 -214
rect -74 -1241 -71 -154
rect -11 -215 -8 -15
rect 301 -215 304 -207
rect 1012 -211 1015 296
rect -11 -218 304 -215
rect 297 -729 300 -726
rect -74 -1244 303 -1241
rect -292 -1258 296 -1254
<< m2contact >>
rect -126 -115 -121 -110
rect -336 -138 -331 -133
rect -157 -140 -152 -135
rect 300 -730 305 -725
<< metal2 >>
rect -379 1464 1021 1467
rect -379 1305 -376 1464
rect 1018 1462 1021 1464
rect 1018 1459 1039 1462
rect 1012 1334 1025 1338
rect 1012 1330 1016 1334
rect 56 1326 1016 1330
rect -603 1302 -349 1305
rect -603 511 -600 1302
rect 56 1195 60 1326
rect 448 1212 1017 1215
rect -646 508 -600 511
rect -571 1182 -348 1186
rect -646 502 -641 508
rect -646 500 -642 502
rect -645 -270 -642 500
rect -571 485 -567 1182
rect 448 1162 451 1212
rect 1014 1208 1017 1212
rect 53 1159 451 1162
rect 511 1159 577 1162
rect -622 481 -567 485
rect -546 1052 -344 1056
rect 53 1056 56 1159
rect -622 -418 -618 481
rect -546 470 -542 1052
rect 519 1045 578 1048
rect 1015 994 1018 1079
rect 52 991 1018 994
rect -604 466 -542 470
rect -527 928 -347 932
rect 52 931 55 991
rect -604 -536 -600 466
rect -527 442 -523 928
rect 525 926 583 929
rect 45 844 1019 847
rect 45 810 48 844
rect -574 438 -523 442
rect -509 804 -328 808
rect -574 -666 -570 438
rect -509 426 -505 804
rect 526 803 585 806
rect 1016 727 1019 844
rect -557 422 -505 426
rect -496 680 -324 684
rect -557 -782 -553 422
rect -496 409 -492 680
rect 41 607 44 679
rect 41 604 1022 607
rect 1019 602 1022 604
rect -542 405 -492 409
rect -472 550 -320 554
rect -542 -903 -538 405
rect -472 381 -468 550
rect 43 470 48 548
rect 43 465 1025 470
rect -513 377 -468 381
rect -452 426 -301 430
rect -513 -1030 -509 377
rect -452 -1180 -448 426
rect 42 402 46 424
rect 42 398 1017 402
rect 1013 348 1017 398
rect -125 -134 -122 -115
rect -331 -135 -122 -134
rect -331 -137 -157 -135
rect -152 -137 -122 -135
rect 286 -290 317 -286
rect 1571 -336 1593 -332
rect 292 -414 312 -410
rect 292 -418 296 -414
rect 273 -541 313 -540
rect 268 -544 313 -541
rect 1544 -650 1598 -646
rect 294 -800 298 -787
rect 294 -804 314 -800
rect 286 -928 314 -924
rect 1564 -971 1622 -967
rect 220 -1057 315 -1054
rect -452 -1184 314 -1180
rect 1575 -1292 1622 -1288
rect 1590 -1364 1624 -1361
<< m3contact >>
rect 1039 1458 1044 1464
rect 1025 1330 1038 1340
rect -349 1301 -344 1306
rect 56 1190 61 1195
rect -348 1182 -343 1187
rect 1013 1203 1018 1208
rect -344 1052 -339 1057
rect 1014 1079 1019 1084
rect -646 -275 -641 -270
rect 51 1051 56 1056
rect -623 -423 -618 -418
rect -347 928 -342 933
rect 51 926 56 931
rect -605 -541 -600 -536
rect -328 804 -323 809
rect 44 805 49 810
rect 1015 721 1023 727
rect -575 -671 -570 -666
rect -324 680 -319 685
rect 40 679 45 684
rect 1019 597 1024 602
rect -558 -787 -553 -782
rect -320 550 -315 555
rect 42 548 49 555
rect 1025 464 1032 471
rect -543 -908 -538 -903
rect -301 426 -296 431
rect -514 -1035 -509 -1030
rect 40 424 48 430
rect 1012 340 1019 348
rect 278 -292 286 -285
rect 291 -424 297 -418
rect 267 -541 273 -535
rect 308 -671 314 -665
rect 293 -787 298 -782
rect 280 -928 286 -922
rect 215 -1057 220 -1052
<< m123contact >>
rect 1016 296 1021 301
rect -288 252 -283 257
rect -334 229 -329 235
rect -50 92 -45 97
rect 568 92 574 98
rect 1157 -352 1162 -347
<< metal3 >>
rect 569 1440 1035 1444
rect -365 1353 99 1356
rect -365 233 -362 1353
rect -344 1301 25 1305
rect -343 1182 15 1186
rect 56 1182 60 1190
rect -339 1052 11 1056
rect -348 928 -347 932
rect -342 928 13 932
rect -323 804 14 808
rect -319 680 12 684
rect -315 550 10 554
rect -296 426 10 430
rect -287 360 10 364
rect -287 257 -283 360
rect -365 230 -334 233
rect -329 230 -328 233
rect 569 98 573 1440
rect -45 92 568 96
rect 1044 -147 1047 281
rect 1044 -150 1161 -147
rect -641 -274 283 -271
rect 280 -285 283 -274
rect 1158 -347 1161 -150
rect -618 -423 291 -419
rect -600 -540 267 -536
rect -570 -670 308 -666
rect -553 -787 293 -783
rect -538 -908 286 -904
rect 282 -922 286 -908
rect -509 -1035 -499 -1031
rect -504 -1053 -500 -1035
rect -504 -1057 215 -1053
use and2  and2_0
timestamp 1700594004
transform 0 -1 2206 1 0 962
box -36 -31 73 27
use decoder  decoder_0
timestamp 1701328861
transform 0 -1 -281 1 0 12
box -229 -7 245 156
use or2  or2_0
timestamp 1700594004
transform 0 -1 -93 1 0 -101
box -13 -17 76 42
use and_ckt  and_ckt_0
timestamp 1701329101
transform 1 0 266 0 1 876
box -262 -516 264 504
use adder_sub  adder_sub_0
timestamp 1701334167
transform 1 0 627 0 1 -469
box -335 -1008 968 262
use comparator_full_ckt  comparator_full_ckt_0
timestamp 1701341286
transform 1 0 2539 0 1 549
box -1531 -756 -340 1381
<< labels >>
rlabel polysilicon -571 74 -569 76 3 S1
rlabel metal1 -570 55 -570 55 3 S0
rlabel metal3 -317 1354 -317 1354 1 vdd!
rlabel metal3 -215 362 -215 362 1 gnd!
rlabel metal3 10 1302 10 1302 1 a0
rlabel metal3 8 1184 8 1184 1 a1
rlabel metal3 -4 1054 -4 1054 1 a2
rlabel metal3 -2 930 -2 930 1 a3
rlabel metal3 -2 805 -2 805 1 b0
rlabel metal3 -3 682 -3 682 1 b1
rlabel metal3 -5 552 -5 552 1 b2
rlabel metal3 -4 427 -4 427 1 b3
rlabel metal2 548 1160 548 1160 1 and0
rlabel metal2 543 1045 543 1045 1 and1
rlabel metal2 543 927 543 927 1 and2
rlabel metal2 554 805 554 805 1 and3
rlabel metal2 1589 -336 1593 -332 7 sum0
rlabel metal2 1594 -650 1598 -646 7 sum1
rlabel metal2 1618 -971 1622 -967 7 sum2
rlabel metal2 1618 -1292 1622 -1288 7 sum3
rlabel metal2 1621 -1364 1624 -1361 7 carry
rlabel polysilicon 2271 1725 2271 1725 1 a_gr_b
rlabel polysilicon 2210 348 2210 348 1 b_gr_a
rlabel polysilicon 2305 1055 2305 1055 1 a_eq_b
<< end >>
