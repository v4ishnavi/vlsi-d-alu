magic
tech scmos
timestamp 1700594004
<< nwell >>
rect -40 -2 -13 23
rect -3 -2 24 23
rect 33 -2 60 23
rect 71 -2 98 23
<< ntransistor >>
rect -28 -16 -26 -12
rect 9 -16 11 -12
rect 45 -16 47 -12
rect 83 -16 85 -12
<< ptransistor >>
rect -28 4 -26 12
rect 9 4 11 12
rect 45 4 47 12
rect 83 4 85 12
<< ndiffusion >>
rect -29 -16 -28 -12
rect -26 -16 9 -12
rect 11 -16 45 -12
rect 47 -16 83 -12
rect 85 -16 86 -12
<< pdiffusion >>
rect -29 8 -28 12
rect -33 4 -28 8
rect -26 8 -21 12
rect -26 4 -25 8
rect 8 8 9 12
rect 4 4 9 8
rect 11 8 16 12
rect 11 4 12 8
rect 44 8 45 12
rect 40 4 45 8
rect 47 8 52 12
rect 47 4 48 8
rect 82 8 83 12
rect 78 4 83 8
rect 85 8 90 12
rect 85 4 86 8
<< ndcontact >>
rect -33 -16 -29 -12
rect 86 -16 90 -12
<< pdcontact >>
rect -33 8 -29 12
rect -25 4 -21 8
rect 4 8 8 12
rect 12 4 16 8
rect 40 8 44 12
rect 48 4 52 8
rect 78 8 82 12
rect 86 4 90 8
<< polysilicon >>
rect -28 12 -26 27
rect 9 12 11 27
rect 45 12 47 27
rect 83 12 85 27
rect -28 -12 -26 4
rect 9 -12 11 4
rect 45 -12 47 4
rect 83 -12 85 4
rect -28 -23 -26 -16
rect 9 -23 11 -16
rect 45 -23 47 -16
rect 83 -23 85 -16
<< polycontact >>
rect -29 27 -25 31
rect 8 27 12 31
rect 44 27 48 31
rect 82 27 86 31
<< metal1 >>
rect -29 31 -25 34
rect 8 31 12 34
rect 44 31 48 34
rect 82 31 86 34
rect -40 20 117 23
rect -32 12 -29 20
rect 5 12 8 20
rect 41 12 44 20
rect 79 12 82 20
rect -25 -5 -22 4
rect 12 -5 15 4
rect 48 -5 51 4
rect 86 -5 89 4
rect -25 -8 116 -5
rect 138 -8 146 -5
rect 87 -12 90 -8
rect -33 -27 -30 -16
rect 111 -25 118 -22
rect 111 -26 114 -25
rect -33 -28 91 -27
rect 110 -28 114 -26
rect -33 -29 114 -28
rect -33 -31 113 -29
rect -33 -32 91 -31
use not  not_0
timestamp 1700473189
transform 1 0 127 0 1 8
box -12 -33 12 15
<< end >>
