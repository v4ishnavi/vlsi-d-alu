magic
tech scmos
timestamp 1700594004
<< nwell >>
rect -5 66 23 87
rect 32 66 60 87
rect 72 63 96 87
rect 125 65 153 86
rect 162 65 190 86
rect 202 62 226 86
rect 249 62 277 83
rect 286 62 314 83
rect 326 59 350 83
<< ntransistor >>
rect 7 51 9 55
rect 44 51 46 55
rect 83 47 85 51
rect 137 50 139 54
rect 174 50 176 54
rect 213 46 215 50
rect 261 47 263 51
rect 298 47 300 51
rect 337 43 339 47
<< ptransistor >>
rect 7 72 9 80
rect 44 72 46 80
rect 83 70 85 78
rect 137 71 139 79
rect 174 71 176 79
rect 213 69 215 77
rect 261 68 263 76
rect 298 68 300 76
rect 337 66 339 74
<< ndiffusion >>
rect 6 51 7 55
rect 9 51 44 55
rect 46 51 47 55
rect 81 47 83 51
rect 85 47 86 51
rect 136 50 137 54
rect 139 50 174 54
rect 176 50 177 54
rect 211 46 213 50
rect 215 46 216 50
rect 260 47 261 51
rect 263 47 298 51
rect 300 47 301 51
rect 335 43 337 47
rect 339 43 340 47
<< pdiffusion >>
rect 6 76 7 80
rect 2 72 7 76
rect 9 76 14 80
rect 9 72 10 76
rect 43 76 44 80
rect 39 72 44 76
rect 46 76 51 80
rect 46 72 47 76
rect 82 74 83 78
rect 78 70 83 74
rect 85 74 86 78
rect 85 70 90 74
rect 136 75 137 79
rect 132 71 137 75
rect 139 75 144 79
rect 139 71 140 75
rect 173 75 174 79
rect 169 71 174 75
rect 176 75 181 79
rect 176 71 177 75
rect 212 73 213 77
rect 208 69 213 73
rect 215 73 216 77
rect 215 69 220 73
rect 260 72 261 76
rect 256 68 261 72
rect 263 72 268 76
rect 263 68 264 72
rect 297 72 298 76
rect 293 68 298 72
rect 300 72 305 76
rect 300 68 301 72
rect 336 70 337 74
rect 332 66 337 70
rect 339 70 340 74
rect 339 66 344 70
<< ndcontact >>
rect 2 51 6 55
rect 47 51 51 55
rect 77 47 81 51
rect 86 47 90 51
rect 132 50 136 54
rect 177 50 181 54
rect 207 46 211 50
rect 216 46 220 50
rect 256 47 260 51
rect 301 47 305 51
rect 331 43 335 47
rect 340 43 344 47
<< pdcontact >>
rect 2 76 6 80
rect 10 72 14 76
rect 39 76 43 80
rect 47 72 51 76
rect 78 74 82 78
rect 86 74 90 78
rect 132 75 136 79
rect 140 71 144 75
rect 169 75 173 79
rect 177 71 181 75
rect 208 73 212 77
rect 216 73 220 77
rect 256 72 260 76
rect 264 68 268 72
rect 293 72 297 76
rect 301 68 305 72
rect 332 70 336 74
rect 340 70 344 74
<< polysilicon >>
rect 7 80 9 90
rect 44 80 46 91
rect 83 78 85 81
rect 137 79 139 89
rect 174 79 176 90
rect -22 36 -20 58
rect 7 55 9 72
rect 44 55 46 72
rect 213 77 215 80
rect 83 58 85 70
rect 79 56 85 58
rect 83 51 85 56
rect 7 47 9 51
rect 44 47 46 51
rect 83 44 85 47
rect 99 34 101 56
rect 137 54 139 71
rect 174 54 176 71
rect 261 76 263 86
rect 298 76 300 87
rect 213 57 215 69
rect 337 74 339 77
rect 209 55 215 57
rect 213 50 215 55
rect 137 46 139 50
rect 174 46 176 50
rect 213 43 215 46
rect 227 34 229 55
rect 261 51 263 68
rect 298 51 300 68
rect 337 54 339 66
rect 333 52 339 54
rect 337 47 339 52
rect 261 43 263 47
rect 298 43 300 47
rect 337 40 339 43
rect 351 30 353 52
<< polycontact >>
rect 6 90 10 94
rect 43 91 47 95
rect 136 89 140 93
rect 173 90 177 94
rect 260 86 264 90
rect 297 87 301 91
rect -24 58 -20 62
rect 75 55 79 59
rect 98 56 102 60
rect 205 54 209 58
rect 226 55 230 59
rect 329 51 333 55
rect 350 52 354 56
<< metal1 >>
rect -118 108 275 112
rect -118 100 -114 108
rect -81 100 -77 102
rect 6 94 10 108
rect 43 95 47 97
rect 136 93 140 108
rect -30 89 -4 90
rect 173 94 177 98
rect 260 90 264 108
rect -30 87 -2 89
rect -30 86 128 87
rect 297 91 301 95
rect -5 85 250 86
rect -5 84 252 85
rect 3 80 6 84
rect 40 80 43 84
rect 79 78 82 84
rect 125 83 252 84
rect 133 79 136 83
rect 170 79 173 83
rect 209 77 212 83
rect 226 82 350 83
rect 249 80 350 82
rect 10 63 13 72
rect 47 63 50 72
rect 10 60 68 63
rect 47 55 50 60
rect 65 59 68 60
rect 86 59 89 74
rect 257 76 260 80
rect 294 76 297 80
rect 140 62 143 71
rect 177 62 180 71
rect 65 55 75 59
rect 86 56 98 59
rect 140 59 198 62
rect 102 56 104 59
rect 86 51 89 56
rect 177 54 180 59
rect 195 58 198 59
rect 216 58 219 73
rect 333 74 336 80
rect 264 59 267 68
rect 301 59 304 68
rect 195 54 205 58
rect 216 55 226 58
rect 230 55 234 58
rect 264 56 322 59
rect 2 45 5 51
rect 216 50 219 55
rect 301 51 304 56
rect 319 55 322 56
rect 340 55 343 70
rect 319 51 329 55
rect 340 52 350 55
rect 354 52 358 55
rect -30 42 70 45
rect 78 42 81 47
rect 132 44 135 50
rect 340 47 343 52
rect 130 42 200 44
rect 67 41 200 42
rect 208 41 211 46
rect 256 41 259 47
rect 67 39 133 41
rect 197 38 324 41
rect 332 38 335 43
rect 321 35 350 38
use and2  and2_0
timestamp 1700594004
transform 1 0 -93 0 1 73
box -36 -31 73 27
<< end >>
